entity uvvm is
end entity uvvm;

architecture rtl of uvvm is

begin

end architecture rtl;
