library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity modmul_control is
end entity modmul_control;

architecture rtl of modmul_control is

begin

end architecture rtl;
