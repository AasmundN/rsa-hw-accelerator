library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity modmul_controlpath is
end entity modmul_controlpath;

architecture rtl of modmul_controlpath is

begin

end architecture rtl;
