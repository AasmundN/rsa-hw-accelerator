library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity rsa_core_datapath is
  port (
    clk   : in    std_logic;
    reset : in    std_logic
  );
end entity rsa_core_datapath;

architecture rtl of rsa_core_datapath is

begin

end architecture rtl;
