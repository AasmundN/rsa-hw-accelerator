library ieee;
use ieee.std_logic_1164.all;

entity foobar is
end entity foobar;

architecture rtl of foobar is
  
begin
  
  
  
end architecture rtl;
